----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:41:18 03/25/2020 
-- Design Name: 
-- Module Name:    FourBitAdder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FourBitAdder is
   Port ( 
		A 		: in  STD_LOGIC_VECTOR (3 downto 0);
      B 		: in  STD_LOGIC_VECTOR (3 downto 0);
		INC 	: in 	STD_LOGIC;
      SUM 	: out  STD_LOGIC_VECTOR (3 downto 0);
	);

end FourBitAdder;

architecture Behavioral of FourBitAdder is

begin

	SUM <= 

end Behavioral;

